module xor_gate(op,a,b);
input a,b;
output op;
assign op=a^b;
endmodule